----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    17:56:21 08/26/2017 
-- Design Name: 
-- Module Name:    ramShip - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ramLose is
    Port ( --clk_i : in  STD_LOGIC;
           addrOUT_i : in  STD_LOGIC_VECTOR (4 downto 0);
           data_o : out  STD_LOGIC_VECTOR (0 to 139));
end ramLose;

architecture Behavioral of ramLose is

	type ram_type is array (22 downto 0) of std_logic_vector (0 to 139);
   signal RAM : ram_type;
	signal dataOUT : STD_LOGIC_VECTOR (0 to 139);

begin
	
	data_o <= dataOUT;
	
	--process (clk_i)
	--begin
		--if (clk_i'event and clk_i = '1') then
			RAM(0) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(1) <= "11110000111100000000111111111111000000001111000011110000000000000000111100000000000000001111111111110000000000111111111110000000111111111111";
			RAM(2) <= "11110000111100000000111111111111000000001111000011110000000000000000111100000000000000001111111111110000000000111111111110000000111111111111";
			RAM(3) <= "11110000111100000000111100001111000000001111000011110000000000000000111100000000000000001111000011110000000011110000000000000000111100000000";
			RAM(4) <= "11110000111100000000111100001111000000001111000011110000000000000000111100000000000000001111000011110000000011110000000000000000111100000000";
			RAM(5) <= "11110000111100000000111100001111000000001111000011110000000000000000111100000000000000001111000011110000000011110000000000000000111100000000";
			RAM(6) <= "11110000111100000000111100001111000000001111000011110000000000000000111100000000000000001111000011110000000011110000000000000000111100000000";
			RAM(7) <= "11110000111100000000111100001111000000001111000011110000000000000000111100000000000000001111000011110000000011110000000000000000111100000000";
			RAM(8) <= "11110000111100000000111100001111000000001111000011110000000000000000111100000000000000001111000011110000000011110000000000000000111100000000";
			RAM(9) <= "11110000111100000000111100001111000000001111000011110000000000000000111100000000000000001111000011110000000011110000000000000000111100000000";
			RAM(10) <= "11110000111100000000111100001111000000001111000011110000000000000000111100000000000000001111000011110000000011110000000000000000111100000000";
			RAM(11) <= "11110000111100000000111100001111000000001111000011110000000000000000111100000000000000001111000011110000000000111111110000000000111111111111";
			RAM(12) <= "00111111110000000000111100001111000000001111000011110000000000000000111100000000000000001111000011110000000000111111110000000000111111111111";
			RAM(13) <= "00111111110000000000111100001111000000001111000011110000000000000000111100000000000000001111000011110000000000000000111100000000111100000000";
			RAM(14) <= "00001111000000000000111100001111000000001111000011110000000000000000111100000000000000001111000011110000000000000000111100000000111100000000";
			RAM(15) <= "00001111000000000000111100001111000000001111000011110000000000000000111100000000000000001111000011110000000000000000111100000000111100000000";
			RAM(16) <= "00001111000000000000111100001111000000001111000011110000000000000000111100000000000000001111000011110000000000000000111100000000111100000000";
			RAM(17) <= "00001111000000000000111100001111000000001111000011110000000000000000111100000000000000001111000011110000000000000000111100000000111100000000";
			RAM(18) <= "00001111000000000000111100001111000000001111000011110000000000000000111100000000000000001111000011110000000000000000111100000000111100000000";
			RAM(19) <= "00001111000000000000111100001111000000001111000011110000000000000000111100000000000000001111000011110000000000000000111100000000111100000000";
			RAM(20) <= "00001111000000000000111100001111000000001111000011110000000000000000111100000000000000001111000011110000000000000000111100000000111100000000";
			RAM(21) <= "00001111000000000000111111111111000000001111111111110000000000000000111111111111000000001111111111110000000111111111110000000000111111111111";
			RAM(22) <= "00001111000000000000111111111111000000001111111111110000000000000000111111111111000000001111111111110000000111111111110000000000111111111111";

			
		--end if;
	--end process;

	-- beres instantno, vrstico ki naslovis z addrOUT_i
	dataOUT <= RAM(conv_integer(addrOUT_i));


end Behavioral;

