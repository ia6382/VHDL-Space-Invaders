----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    17:56:21 08/26/2017 
-- Design Name: 
-- Module Name:    ramShip - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ramShield is
    Port ( --clk_i : in  STD_LOGIC;
           addrOUT_i : in  STD_LOGIC_VECTOR (5 downto 0);
           data_o : out  STD_LOGIC_VECTOR (0 to 74));
end ramShield;

architecture Behavioral of ramShield is

	type ram_type is array (47 downto 0) of std_logic_vector (0 to 74);
   signal RAM : ram_type;
	signal dataOUT : STD_LOGIC_VECTOR (0 to 74);

begin
	
	data_o <= dataOUT;
	
	--process (clk_i)
	--begin
		--if (clk_i'event and clk_i = '1') then
			RAM(0) <= "000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(1) <= "000011111111111111111111111111111111111111111111111111111111111111111110000";
			RAM(2) <= "000011111111111111111111111111111111111111111111111111111111111111111110000";
			RAM(3) <= "001111111111111111111111111111111111111111111111111111111111111111111111100";
			RAM(4) <= "001111111111111111111111111111111111111111111111111111111111111111111111100";
			RAM(5) <= "111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(6) <= "111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(7) <= "111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(8) <= "111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(9) <= "111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(10) <= "111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(11) <= "111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(12) <= "111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(13) <= "111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(14) <= "111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(15) <= "111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(16) <= "111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(17) <= "111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(18) <= "111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(19) <= "111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(20) <= "111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(21) <= "111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(22) <= "111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(23) <= "111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(24) <= "111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(25) <= "111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(26) <= "111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(27) <= "111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(28) <= "111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(29) <= "111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(30) <= "111111111111111111111111111111111111111111111111111111111111111111111111111";
			RAM(31) <= "111111111111111111111111111100000000000000000011111111111111111111111111111";
			RAM(32) <= "111111111111111111111111111100000000000000000011111111111111111111111111111";
			RAM(33) <= "111111111111111111111111110000000000000000000000111111111111111111111111111";
			RAM(34) <= "111111111111111111111111110000000000000000000000111111111111111111111111111";
			RAM(35) <= "111111111111111111111111000000000000000000000000001111111111111111111111111";
			RAM(36) <= "111111111111111111111111000000000000000000000000001111111111111111111111111";
			RAM(37) <= "111111111111111111111111000000000000000000000000001111111111111111111111111";
			RAM(38) <= "111111111111111111111111000000000000000000000000001111111111111111111111111";
			RAM(39) <= "111111111111111111111111000000000000000000000000001111111111111111111111111";
			RAM(40) <= "111111111111111111111111000000000000000000000000001111111111111111111111111";
			RAM(41) <= "111111111111111111111111000000000000000000000000001111111111111111111111111";
			RAM(42) <= "111111111111111111111111000000000000000000000000001111111111111111111111111";
			RAM(43) <= "111111111111111111111111000000000000000000000000001111111111111111111111111";
			RAM(44) <= "111111111111111111111111000000000000000000000000001111111111111111111111111";
			RAM(45) <= "111111111111111111111111000000000000000000000000001111111111111111111111111";
			RAM(46) <= "111111111111111111111111000000000000000000000000001111111111111111111111111";
			RAM(47) <= "111111111111111111111111000000000000000000000000001111111111111111111111111";
			
		--end if;
	--end process;

	-- beres instantno, vrstico ki naslovis z addrOUT_i
	dataOUT <= RAM(conv_integer(addrOUT_i));


end Behavioral;

