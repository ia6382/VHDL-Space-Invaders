----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    17:56:21 08/26/2017 
-- Design Name: 
-- Module Name:    ramShip - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ramWin is
    Port ( --clk_i : in  STD_LOGIC;
           addrOUT_i : in  STD_LOGIC_VECTOR (4 downto 0);
           data_o : out  STD_LOGIC_VECTOR (0 to 62));
end ramWin;

architecture Behavioral of ramWin is

	type ram_type is array (22 downto 0) of std_logic_vector (0 to 62);
   signal RAM : ram_type;
	signal dataOUT : STD_LOGIC_VECTOR (0 to 62);

begin
	
	data_o <= dataOUT;
	
	--process (clk_i)
	--begin
		--if (clk_i'event and clk_i = '1') then
			RAM(0) <= "000000000000000000000000000000000000000000000000000000000000000";
			RAM(1) <= "111100000000000011110000000011110000000011110000000000000001111";
			RAM(2) <= "111100000000000011110000000011110000000011110000000000000001111";
			RAM(3) <= "111100000000000011110000000011110000000011110000000000000001111";
			RAM(4) <= "111100000000000011110000000011110000000011110000000000000001111";
			RAM(5) <= "111100001111000011110000000011110000000011111111000000000001111";
			RAM(6) <= "111100001111000011110000000011110000000011111111000000000001111";
			RAM(7) <= "111100001111000011110000000011110000000011110011110000000001111";
			RAM(8) <= "111100001111000011110000000011110000000011110011110000000001111";
			RAM(9) <= "111100001111000011110000000011110000000011110000111100000001111";
			RAM(10) <= "111100001111000011110000000011110000000011110000111100000001111";
			RAM(11) <= "111100001111000011110000000011110000000011110000011110000001111";
			RAM(12) <= "111100001111000011110000000011110000000011110000011110000001111";
			RAM(13) <= "111100001111000011110000000011110000000011110000000111100001111";
			RAM(14) <= "111100001111000011110000000011110000000011110000000111100001111";
			RAM(15) <= "111100001111000011110000000011110000000011110000000001111001111";
			RAM(16) <= "111100001111000011110000000011110000000011110000000001111001111";
			RAM(17) <= "111100001111000011110000000011110000000011110000000000011111111";
			RAM(18) <= "111100001111000011110000000011110000000011110000000000011111111";
			RAM(19) <= "111100001111000011110000000011110000000011110000000000000001111";
			RAM(20) <= "111100001111000011110000000011110000000011110000000000000001111";
			RAM(21) <= "111111111111111111110000000011110000000011110000000000000001111";
			RAM(22) <= "111111111111111111110000000011110000000011110000000000000001111";

			
		--end if;
	--end process;

	-- beres instantno, vrstico ki naslovis z addrOUT_i
	dataOUT <= RAM(conv_integer(addrOUT_i));


end Behavioral;

